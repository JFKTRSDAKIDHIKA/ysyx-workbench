module bitrev (
  input  sck,
  input  ss,
  input  mosi,
  output reg miso
);

  // Internal signal declaration
  localparam IDLE = 2'b00,
             RX   = 2'b01,
             TX   = 2'b10;
  reg [7:0]  counter;
  reg [7:0]  data_in;
  reg [1:0]  state;
  wire inactive = ss;

  always @(posedge sck or ss) begin
    if (inactive) begin 
      // $write("inactive\n");
      state <= RX;
      counter <= 8'd0;
      data_in <= 8'd0;
    end else begin
      $write("active\n");
      case (state)
        IDLE:  begin
          miso <= 1'b1;  // slave空闲时, 将MISO信号设置为高电平
          state <= IDLE;
          counter <= 8'd0;
          $write("IDLE");
        end
        RX: begin
          $write("RX");
          data_in <= { data_in[6:0], mosi };
          counter <= (counter < 8'd7 ) ? counter + 8'd1 : 8'd0;
          state <= (counter == 8'd7 ) ? TX : state;
          miso <= 1'b1;
        end
        TX: begin
          $write("TX");
          counter <= (counter < 8'd7 ) ? counter + 8'd1 : 8'd0;
          state <= (counter == 8'd7 ) ? IDLE : state;
          miso <= data_in[7];
          data_in <= {data_in[6:0], 1'b0};
        end 
        default: begin
          state <= state;
          $write("Invalid state");
          $fatal;
        end
      endcase
    end
  end

endmodule
